`include "Defines.v"
module memory_control (
    
);
    
endmodule